module memory(

input save,

input[3:0] save0,
input[3:0] save1,
input[3:0] save2,
input[3:0] save3,
input[3:0] save4,
input[3:0] save5,
input[3:0] save6,

output[3:0] number0,
output[3:0] number1,
output[3:0] number2,
output[3:0] number3

);


endmodule
